library verilog;
use verilog.vl_types.all;
entity \register\ is
    port(
        rs              : in     vl_logic_vector(4 downto 0);
        rt              : in     vl_logic_vector(4 downto 0);
        rd              : in     vl_logic_vector(4 downto 0);
        writedata       : in     vl_logic_vector(31 downto 0);
        regwrite        : in     vl_logic;
        A               : out    vl_logic_vector(31 downto 0);
        B               : out    vl_logic_vector(31 downto 0)
    );
end \register\;
