library verilog;
use verilog.vl_types.all;
entity test_alucontrol is
end test_alucontrol;
