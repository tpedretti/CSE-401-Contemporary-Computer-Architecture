library verilog;
use verilog.vl_types.all;
entity mem_test is
end mem_test;
