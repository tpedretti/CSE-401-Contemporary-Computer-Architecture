library verilog;
use verilog.vl_types.all;
entity adder is
    port(
        add_in1         : in     vl_logic_vector(31 downto 0);
        add_in2         : in     vl_logic_vector(31 downto 0);
        add_out         : out    vl_logic_vector(31 downto 0)
    );
end adder;
