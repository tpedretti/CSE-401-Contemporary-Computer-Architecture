library verilog;
use verilog.vl_types.all;
entity test_mux is
end test_mux;
