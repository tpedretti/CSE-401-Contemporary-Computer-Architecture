library verilog;
use verilog.vl_types.all;
entity idecode_tb is
end idecode_tb;
