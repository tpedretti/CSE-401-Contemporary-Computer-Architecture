library verilog;
use verilog.vl_types.all;
entity pipeline is
end pipeline;
